module main

import hall_of_code.vping

fn main()
{
	println(vping.ping(ip: "hosting.ottnec.de"))
}